`timescale 1ns / 1ps  // ָ�������ʱ�䵥λΪ1���룬ʱ�侫��Ϊ1Ƥ�롣

// ����ģ��dff����ģ������ʵ��һ��4λ���D������
module dff(
    output reg [3:0] q,  // ����˿�q��4λ�Ĵ������洢�������ĵ�ǰ״̬
    input [3:0] d,       // ����˿�d��4λ���������ô�������Ŀ��״̬
    input clk,           // ����ʱ���ź�clk������ͬ��״̬����
    input rst,           // ���븴λ�ź�rst���������ô�����״̬����ʼֵ
    input en             // ����ʹ���ź�en�������Ƿ���´�������״̬
);

// ��������������Ϊ��always����ʱ���ź�clk�������ش���
always @(posedge clk) begin
    if (rst) 
        q <= 4'b0001;       // �����λ�źż�������q����Ϊ0001
    else if (en) 
        q <= d;             // ���ʹ���źż��������d��ֵ�������q
end

endmodule
