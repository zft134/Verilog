`timescale 1ns / 1ps  // ����ʱ�䵥λΪ1���룬ʱ�侫��Ϊ1Ƥ�룬���ڷ��滷����

module FSMTestbench;  // ����ģ��FSMTestbench������һ������ƽ̨ģ�顣

reg x, y, rst, clk;  // ��������Ĵ�����ʱ���ź�
wire z;  // ���������

FSM fsm(  // ʵ��������״̬��FSM�������Ӷ˿�
    .x(x),  // ����˿�x
    .y(y),  // ����˿�y
    .z(z),  // ����˿�z
    .clk(clk)  // ʱ���ź�
);

initial clk = 0;  // ��ʼ��ʱ���ź�Ϊ0
always #5 clk = ~clk;  // ÿ5��ʱ�䵥λʱ���ź�ȡ��һ��

// ��������
initial begin
    #10 rst = 1; x = 0; y = 0;  // 10��ʱ�䵥λ�����ø�λ�ź�Ϊ1��x��yΪ0
    #10 rst = 0;  // 10��ʱ�䵥λ��ȡ����λ�ź�

    // ��ͬ������벢�۲����״̬�仯
    #10 x = 1; y = 0;  // 10��ʱ�䵥λ������xΪ1��yΪ0
    #10 x = 1; y = 0;  // 10��ʱ�䵥λ���ٴ�����xΪ1��yΪ0
    #10 x = 0; y = 1;  // 10��ʱ�䵥λ������xΪ0��yΪ1
    #10 x = 0; y = 1;  // 10��ʱ�䵥λ���ٴ�����xΪ0��yΪ1

    #10 rst = 1; x = 0; y = 0;  // 10��ʱ�䵥λ���������ø�λ�ź�Ϊ1��x��yΪ0
    #10 rst = 0;  // 10��ʱ�䵥λ��ȡ����λ�ź�
    #10 x = 0; y = 1;  // 10��ʱ�䵥λ������xΪ0��yΪ1
    #10 x = 1; y = 0;  // 10��ʱ�䵥λ������xΪ1��yΪ0
    #10 x = 1; y = 0;  // 10��ʱ�䵥λ���ٴ�����xΪ1��yΪ0
    #10 x = 0; y = 1;  // 10��ʱ�䵥λ���ٴ�����xΪ0��yΪ1

    $stop;  // ֹͣ����
end

// ����������ڲ�״̬
initial begin
    $monitor("Time=%t, rst=%b, x=%b, y=%b, z=%b, state=%b", $time, rst, x, y, z, fsm.state);
    // ʹ��$monitor���ٺ���ʾʱ�䣬��λ�źţ�����x, y�����z�Լ�״̬����ǰ״̬
end

endmodule
